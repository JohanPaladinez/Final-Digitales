library verilog;
use verilog.vl_types.all;
entity Cod9a4 is
    port(
        A0              : out    vl_logic;
        N1              : in     vl_logic;
        N5              : in     vl_logic;
        N3              : in     vl_logic;
        N7              : in     vl_logic;
        N9              : in     vl_logic;
        A1              : out    vl_logic;
        N6              : in     vl_logic;
        N2              : in     vl_logic;
        A2              : out    vl_logic;
        N4              : in     vl_logic;
        A3              : out    vl_logic;
        N8              : in     vl_logic;
        M               : out    vl_logic;
        N0              : in     vl_logic
    );
end Cod9a4;
