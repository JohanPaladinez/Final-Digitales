library verilog;
use verilog.vl_types.all;
entity Maquina_estado_vlg_check_tst is
    port(
        W0              : in     vl_logic;
        W1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Maquina_estado_vlg_check_tst;
