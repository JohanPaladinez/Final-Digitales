library verilog;
use verilog.vl_types.all;
entity Nuevo_4a2_vlg_check_tst is
    port(
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Nuevo_4a2_vlg_check_tst;
