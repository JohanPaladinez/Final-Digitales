library verilog;
use verilog.vl_types.all;
entity Nuevo_4a2_vlg_vec_tst is
end Nuevo_4a2_vlg_vec_tst;
