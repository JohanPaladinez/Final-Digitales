library verilog;
use verilog.vl_types.all;
entity Comparador_vlg_check_tst is
    port(
        D0              : in     vl_logic;
        U0              : in     vl_logic;
        U1              : in     vl_logic;
        U2              : in     vl_logic;
        U3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Comparador_vlg_check_tst;
