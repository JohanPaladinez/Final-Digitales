library verilog;
use verilog.vl_types.all;
entity Cod9a4_vlg_vec_tst is
end Cod9a4_vlg_vec_tst;
