library verilog;
use verilog.vl_types.all;
entity Nuevo_4a2 is
    port(
        Y1              : out    vl_logic;
        F3              : in     vl_logic;
        F1              : in     vl_logic;
        Y2              : out    vl_logic;
        F2              : in     vl_logic;
        F0              : in     vl_logic
    );
end Nuevo_4a2;
